��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]���9w��VpL���~�����.��7
���l�g�S��N.���c����`��8��:��!�o�L�����P�Z�:\��P�&z-���,¾��DF�@��IJ:O�B$���nG��fx`x}�����N&�5b̸�Z�*���ʄ����	߈�R�6�N��+! �ch���c�qb�!��,��2P�2�W1j9��n���C�A�05�l����cn��Ɩ�Ur �coGͰ�ء�9�	�ӓ���&2 ����d/�*Q&T���	�@d�҇j�
�w���/����s�/p�,<�;�'�i�ϸj�\og̓(��X�>��y���~3�[Q*fA��m_�X�0��ϑR�.���Efg.�s
�
_FrA�C�&�A��l�u�mm�%�T�v�|o?,���y���s�!+�-�k���.f�<.�PE �lr\�����B��pW���3��
~��;4���湂���
Ռ���č�]��[���"v2�2q�^T���7�-	�8�ƤS,�ʡW9���J�p�)IR�� G�&�D��"�K�2g�j8	H��Mڍ�0�
���j@N��=����>MIˇs�=y�����hy�leGgp'~�L�MSh�`�>E���|�_��\��N��0V�=�{+*7I�,+l~������.��5מ]t��uj��z�|?i����;����D������N�����73���n�~�����:X��%�����Xf�/�&���~Q�i�C���e�}B�7N������$P�Jk��i�8����%$wRc �Tp!?�e�c{H�rC��������]GM�7�kk�������l�v��F#oWt#�y�>������V⸰f<��ޕFd˟�!2�.�IT����$ ����>�W/@\	J:��T;���|�	�H+I��nGWQ֌$�<�� >0�>��A�C����KL-���fT���������o̢��.h��;	�3��	���'9$H-�~�#F ����0Vb)IIL�R<d��F��yV����7W�����"�qS�o�[�S�K��&���H�껫���1.���I��Y�[�,�:Y��*5�tq�9��hj3�IB�����~�S���O/t����Y����O���m���n%b���e��ě=�rN�`=b��}/Ma�)�f��&��ߪj0��cL9��U��2k'�^�N���vr�M�����j �F�b��V�ba|�m�	�+��E$i��:z�bXI5Mb-�}���ك��j�wШ��Y��|Fr��!/���a��A:�>�������m����]L��«��r�M��a�X5"��[��h�y�k�Qx-l9�b6t�J@&�Ҍ�%�]�����]�9������9N8��B|��{c�E���u
�C�@�8�U��3�.?٨��h#�m�Ǧ���Y�,+k�k��럝$����
�I	�R>�JَߺƟ�n;�}�3Y��,�ϻ�����7��Åǩ��n�8{��I�G0C�`�dAE�ٗ6F_�Qc��Ne����:g�m���<=o��MW(m����m����<�2��dZ����؛I�*5Q�]�m�ު�v��>�(;	�F�[�@��~3R���:�P�]�ѱ:�����6/�x��&F8ٱww��T��y���1����'m�Ѽ.$
��|��=_c:��L�~��u���2�֟b�E83	��ւ�Qܷ+v�_�ʅ���ވ�ݾ��l@�� ��.M�aKŘ�F>�7/�x�:��V��X|���TW��̸���kk�)*�̏�G\�v��f`��s(��|��C���,�COH����1@{{�d�2�rU����y>�I��.o x��گh/����u/�W6#h^�"7���k���4)>���¶;꥜]VBѯ�in��z�*8"Gv��C��(n�<wNP��^�$^
=f���'
ƀ�j�HU��$�����8�P{FA̦G�Ů�`�2.����?/!���^_�Ű��]�=��7x�?����!�Lcf��b���:5����JX��1�М���S�R��ܺ��:�ncU8^��6��诹�ɂ�l>����*�EX�*
f�vQI�!:^#����w��-�b����G�-%��������؟[��Ȗļ?�Vn۲C�4un��0G2��']u���>�)�K����<2��@ޙ_C�7㷨�N��R�NL��#����l�&��vjx��ޛ�H5�>�b�l�Y(I�l0�.�|�\!�;���>���^�(l�>fb�[�V����5̴;l\�?�f����ȿ�}���t1Q�kbջ��Zk�`)�Pv31���B�Jb �eW�;�l9�����M_���!4�_P���B{|"n� p�p�e��{0��Ԫ�)��&`��
�?D�-�l"ȉ��tƾ��T�,�^�>��&�c��@q���cHecÚ�^���[��״�䰄������EAʈ�	ϸ��T�r��Vzw��q���'UL���iMб��̇����O�T1X�A?�Q�k@�Hw��vX�����Bm_�yq݁o��FvqĦ��[N�*,f�[���2?�65�\�JY=!���4Jr'�@WR�cq��0�q8��
�1^�����\<�[�����d��I;mǠ�<*$����/�p0.��^NY:H5� ���r9�ڳ<�Ɩo"19(M>S>W"�&���qK�M���^�M�Q x8��@u�h�[|1]�C�U�D{2%�H_��,���>C�:���F->9�E0=W�;��ٽ��ڝ˪���,a��VlH��h�=ܥu��V����w��?��`T��H�wE$�W�����֒����$��v�}aRl�M ��naZ�W�v�=C��_���_'��C!����s�Aa�B�e5�o6�C����f��s�//�=c�|�`�����n4:�������1�%�쟋m�B�}�=��Ǚg���N��Fq��ġ�B��	�C6���/���A�ʏ�����\b� ���+�`�����頂x��TrޣW[dy��r�L�cL���!d�M�r����i ����[ס��v���ȃ����R���B���`B<�_��4�Y۹�ZX2l�bB�\�k�w7lD6K0˶��gZ�vI��9��2�5nΔ_I�,��nI"�t�>���q��]^S&���sc�L �+��}1cF�R�?#�~��Ex��&�mkl��_�]`�栄k��4����_��5xL���s;!�}|q�_z�?���g����Gx�	M�Į��Q����c�g6\�VA�]�yT���l�����G�A����M�g~Tx~��cUG^�JVF�m�am����!�Ѣ�x�n�d��	H���!�Z���A+t�q�? 윎�Y�TW����$��1� ������~��`hbn�L��8��#{���^$��±��U�Ũ�{J/]d4��}Q��[��@�ؾ�u�eUV�_ƽy�����
.� 7Yho��s8O	��'q`���O��X�=�"�ly7�I�Y!)x�,Ak�	~��n�!�=�S�eBn��T��{�)���QD�zA:}�f��-u��2.�`q�S�y�=f����ç��A�)��8�l�|��a*
�w}<����sbW(�E��s2`�'hw0��*��C�K��A���~�@p��"&�8XA��|<S$������}W�&��>,��a����z�\����+�sq�c�g n��uC���6��Ei�ۗ(*�0�F+��,�+Q���c����	M�VF�0��h��H�~J}R���r]S�MC-�8�]�X��=�g�$g=d����'��̈́��/�8q�J���������iK��}F�<��>�/qT���I
���xK�E�������SriB����r���:r�}m.۞�#�e�7�&j��x�)V��Bk�:PNOG�ks��6_�D�QP��.j=I�u��x��!d:���u�0⤟�e/܄��B}U��~]H"~�=�	����fZ��Y2r�:���b��Q�8�S�F��b�YF|��P���b�s-�Äх'J�����[`��]4��W��p�(�d�i��آ�{1l]X����Jq�)�m��"���_-��jQ��|T�u!�us`�X^��Ѹע1S欑jŒr�2&H�(!-H���Yѱ�[w9���n��ϱۚ,C��,Vh38����޹q���'׶+��x�?z�NӑD�B�[���{DUX~�/NWkg�-��{���їWC��L�=r���񶑽Q�	��>2�ܙR�T|�^J��S�p��go��}�Gȿ����Q�+�Z���itJ?�p�)���	;�B�r�˞�o� ��[G9Ȼ���=7;x�Z�g�/5��:��?���$�DX��PK�h����/�`�x�	,J����G?�TR��ݎ�����9����,����4��a�]6���r�<Y��Q?�l��`R���&ѥ�w���`;T?��;	tl<{���ã��R!$D2�1ɲtOs�yx.D���+Ѳ	�hgQs ����V�똶�;B�J,c�DfYZ�3 K�U�z�*l�yjo��K�%#Z��,��ti�$.�ʺZD[�����o�)����4K^Q$~[Q�y��g,��E�d�cX!>[�m޷F��׸s�9I�r�����:�b�O{�9�-MLD?�%"�����W�4��� 3�.�9(N�����1��]-5�"��[/Sa]m����Nأ�".���F��P)��}D����Ut�c��3��Wg�:@�!�5L���E��z^�0W��W.;�"��#�W��,<Dm���-�H��.��M���.<�j$��i�=O�s��B��ǀ��}��t\Xy��.~�f�4�/���:���� ��b_:�p>�wh���Yh7�Aۡ�'��g�����3d,J
�l�2ϕTdZ@��=�@��?J�� Z�R�e��y�U3hC���:�؇&�*Z
��!�2�^_̺���w*f�����t��
��*}&1��6��EJ!�WM[0���xI~E3����fNa�q����8����A/��݈����`ڬ6�E�k��q��'-� ��*�1�n@p$&C��u�	�Gh2�7:х;��`�H���T��6!� �r϶���rhH08��)���2:�-E��,,%���j�,m�7@	���Y�Q�s?��M�H2>ɢ��b�gĐ���ך�Ɨ�ħĀ+�g%b�"����k��tt@���)�.GͣcK2��Yud;�x��+趦��>T��r������"��O��4�߯��
$H]��/���9�ذ�aVkv�[��(5��R;�kTI�Ϧ*W��F&D�6�o ������eɵ�atg:�,4��T��{�S��p��R��|_-�B+������d'좓�ƫӑa��T�v���P���0k�s�$��Q�I��+�����Y��~Xp�}d�l�[��b��%�'�q=��J�OS���0��QG����x-���VS��n7ËOR�s�'�$s�[�k�ՔE�r5���kO��sW6ğ��j#�����Ƣm���*(m��s�[��ԣM�����0=aW����;k����6��y��R�I��x�Ԓ�iAs����ز��� �8?�~�h���Tʠ��V�lf��H���$b�/�,������Q����p�m �
\ʌ���x^T����B����y&%.��U�mw��b��|�5N��vӾ�&Lv%©�HY;����9^����H9�/�U����,6
��py�3��)No1��,�X�Ak�e����%�8u�k ����S�P�Hx�,Q�>ƕ������˶+l�f�Y+0�>VW�3S�s��
���u��N�1���9��1�3I'���o^��[}��A
H5o���!�b3fm�����)^ɤA!�UU��Z�J���t`���:���A�����N��>���pU�ٗ�*�}��2�;o�L�A�R��ү5No�N�#�@���[�;ktP����83ߓɑ�`� 	br=�?��>���p��)�<XV��1q�k���'��ز{��Z]�9�b˲ḅ�^������6/�C&XL$�$�a%� Q��u�s-��(�Z��J�'�tf�0�r��D�Z� a*6�5y�bk����p��jM��jad&�Y��q:)^_Wԟ������C
��!ӽ��uPal:!d
�#R|���ɉ��]�ɸ���A��_�a&0�9�*�R�Fڇ�x	�W.i�:��Xm�xｨ�.��[�ڡ��+K6º�!Lj��t-,�_��DnV"cj��!�Ş�_�3�"�j�����:&��O�?�r�#�eIY����J"tf'���v�"95��Im��yB@��6��S%��Z֏�Bei�N����=~��z(y��x�.�d�>����/��=#{��3�-%*DE��k�Bqd�"<��2� �U��'Jǧ#����W�Ѓ�F���'g%�r���qp�[Ub���*`FFK#�cw���;VV��p׭İ"�R���-;@���¿�k��o�?��������$�k5��^����M�ɮP�r�P@�Pu��������M�&�SsZ�P�R����>Ӥc�3,�%�8�8�ت9�>ٓ��Q��{�&�BXRPՌ�D>��� �� �>2g�v��	ꖿH��{��Q�`�ʂuG���)T3�s���HG�a�!߉�+���D� ���7Ⱥ�*n�Q��.]t�b�c>��0�v	}�=<=�<�n�r�����Ρ߆�R���u�e�1`�m_�g/�Wr��:��~L]b����	�K���Z��.3��0��l�0t&�W�y�B?�1~���G\�A��ɹd���O��i���'�O��&F��Kъ��vr�����\ޘd>^��xU��	�b�8�f��c)rK��c��R�^%�i��:�A$a͉�� t�:ԑ�yd��1	H��{T�\����%U�	��)���B%5׋
�b�@��_F�r�m�`�pb�}��pp	�E,+���-fA6��&2���V�u[C1઴XT$6�I>�[k~Y��X�:��s����+s_NW.8(��}j�]V�Cq�d݉���i�
���,��~1�M>EȦ~�X��]�P }��j����3-:��2��/q�s���%Vf;���v��X�/D(d���O������S3p�1Zc?�L̴&,Y��P4!��u�H��2\��l�M̎�U�O
���v�a��1�����ǹj�{����B�o�k"v���T5tgl�H����)�]0{0��/T:וs�p='B*��e�aQi5B��`Hy�]"����d W��b�̠��2\�n����l�k��f�L��k�J�[�NԶ"3'v��f��߬]ID$�_�O��E���?�o��ZD~�ek��Yԯnv�l��L�Ĵ����g�������{��ƹ�����[ۓ)��[٠�� X=�A��	��h\�����)�!O�  ׅo}az�T	�Xaw����~�8�ׇ�ݼ��#;�03��>��d� ��D>A��:S��,-m��,�����,@)�r���W��m��l�uL��������o3��"���������N�g��^�r�kk�Sޜ�*��Vbbf�K��C�(`qL�Į�������<-툋�6�V��M�u���)������4��!��}�A��e���ν�^����z����?#aj��c4cO7�'�#�_�u�Lގ��+N/���C]ooI=�W�d7�\Ƣ�J���"�av�Q��|��"�wĈ"�)"3/����>�ي������1U�\��-�b_\6�7���� ?r��U30���(������,J�6����=��w����p3ަ�O����Y��9	Nλ�D��
r�<�_�ȝ�8m�(�bZ 񐿃�qwF���������k�~)_��d	��<{d#v�����Eb��)�P]�	χ*�\X��6��'^IZ�E��1�^���h4�6����5r�U��	�W���tғj{/�k��3��{c#����.I8��-v7㴛4A��B�3��4"��mK�rY�4�����u��հ.�U���뗯�VO�E����4��eJ�P��Fw�o���O��_�f�f�~���˵S�r�?����y)��o6����~)�\sBp|�������2�ح&F����v$	I�d�1~�ܠ�H$R���.U�"��>;�ӻ	�2r�4wz����z�� ����vpӟ\��p#]H��`����fϝYg����e��p(�y��"+�('#�^sLa� ��@!eѳ��]�Ԉ)��4[����0f=c��$����%��Z�6�ױup������q$"[���b:K?�I�dh!E0'�)%��^�
>���� z��T�4���
'0��C.�1JV}NU�'<U	*[܅#XBO>�e)+X���Q��l#�n�ң��ɗ�o]sZ��ҍ�_�0Z2W8���m=��g/�H<jr��;Ih`yP�B�Q��x�I����	T� "�c.K�"��f�t�.<2��\��)�׏5κ!=�E(A�l�փ���NS�5>r�4o��"/��"M�J��#���$U��F���G��\���Ω�|�u��gA�/��E�T�dC��W�J�:��@W)�G��"��P{k�0?�7��T���z�&�\�CP�(�İ��8Cz.�]�nb�V��!�̫-<�Iu"`�Cʪ���Nk�VH�Y���:��$.ᗡ���xʋ����h�5��y<Cڇ���h^Sxy{�Ϯ�qD�Y�����ib␠�Q�,t�`��[�`%�V��6�؞,_���S�}W�"�ڵ��3�ϻ��P��4��t���֌;ͯpI���k�A�TF�e�DJ\S��/	9I�c�j@�P8�!`V��x��b��1��!��G���U��+�>��|�d��%φ���l���aPf�Sa��������0�c�n{��E�Z�U7��w� {��������w�����a�c�D�\~w�M��킴9�`Oa��:
r���`4BFI9&�t�G����b�Qt}bc�Yu���o�:f�?]�gV�P',�}ж��)�֔��]��XM炦���D�g]����EgĩZDɏ�-禜���ν��ğhK��cdsr�A���1��[��E�F c�F#!N7>�
�v��j~��f�8"�I�m�y~�w$�2�}�n�⩅�#3���5?{��$�8*]1�_M`�;�j�bXq���Lx2D��[)��2H ����Z�l�7ȹ���h !t���wC�����D(�Ngp���45�������'�Q�R�jO��n�H{+qf�7�n�|���c(�Fk��Tsm
�)���rͤAaQ=�`sˎ�LW���h3�/�2\����#���T���T¼�O��Q�H�;����ȏ8�����y�2��-��bW��z�;��6q#��Ђs|���.��@4o����=��_�ם�����C��I��D=o��'�k�:u���@��D�,:^o�
�A[8'�"���� 1�c�O�����O  ���W`�I�phn�-��lu����������s��<�`�������*���4��=,K���L��%��5��sx��"P���Qt��%{"ᬧ��8D<��Q��/�E��rB�^|,|g(E���� 3�_�}�{f�c�I�f��������t�՜�YmυL�#��>��/���k����^��e����������j��-J������.��>���A��വ�F��Q�����lo<���A�-2��U�U=����,�������e���B;��C������E��l�����%��%E}���z��Wg���,�@��C3"�P��X�FU��#�&r	�?�SN�N��&��Zm[k�W#�_�闦�eT���ã��.tG�$�8�Pج�h�d�5�3���]t��C�8��+��
�B�k$Tx{�'�Y [0^v*��n�}�6��t瀾8����%�ْ����y����<l��I��Т��Γ���F���e���I�>)-����BӸ��O�@����cV�/L�#|．@x9z'f��O[�ʒu@͕�����B�4�;1����%B����3Q绩��!��~ĕZ�z��kx�f;immٙ�_*z�Z�z�m���@����ae=�:���r� ���'RP�vhۧ(�LǊd�����6M6.�~CQ�� :c4@�.a�s렌`c����mOv����RLz�)�g_��*9�[��n�.��󥷖���(>�V���BP�0���:F��m^R-�0Q����[[b�ړ�^ÞAf~M��2�Q��Q�U(S�7��)�:����DTIZv���g.(=�����X���F�5.�	�O�2�_���k0@sCy���z:�f᫉i�iV���jo�m�$�Z �3wf�!��q�`��v�������S>Z�N��t�mOs����������A�׮~��ܡw����޲�� �~F1���}E'��%��Xt�&ƞ�1;�;�+O��?)� �{+`��4� =1*T�;X��b���N�ֳ 9�z6xE店�o#/�fk}{T�lA���8龰���ێ#�O$���.M���Y��]�u=0����MS^v��2��\�������W��퀡���>��]y���B��E^�yh���fDT�Ȉ56�6X#������(�W<�
y��P����2��քgZ��#Y�l�.^���	��+��*��1��LZ:?����yD����P^�C��I�-��w�ek���U�������TU���M�҉O�"i�*�Ĝ!kW�u6u��KY� �ï�<x>(&�a����.�q��1[����$m�~�ڪ�e� ��m ���y�U�=�����|ԨY*�ȢI����-t*B���`.�S��H����}{�v[1� ��"���=�;�Q�Ȱ?�����i5y6��W����1���Y���*{��gVV"��aOI�����>�rH[G+].�{q��L{��x(��B��7�u���N� ���Mr��J��M��;�
�#����$XNo759;��4�𮵒�q�y�;��P,^��'�4�q�~֎t��ƅ����M6�y&�}v)���D5.���hXP�xoi�Y��a�udS涣/(�®���x�˔�!�.��у��y�r1�ߑG*��X����E���5�AJ����K���z�J(E�?��{��i�Ff��vH��'A��+z%~,XZW T��Z�vۛ���K�d|*;3Ɩޒ7�i���>��%����/��B߅�=߰�����l��V�%�Zs� ��p��P*���D?}FL4�wp��/���'�t�DP�78��𒅪^,qv���<;�M0`�.ߍ_�ic��D�;�4I9	ߕ�F�Zv��ږ��O�q��Wޯ���S>�&���r��J�v�:��d�Q����p�5�X��"Q��f�)+y-G���kCE�E&6P�q=w++���1���G%��@q�<1a|D�T��]��0jv?|�Я8�����&�S�P�s��B�pbR
B�1�	��R���!�-����x�3��D�d�"*��Ű����/�A�IL��kb�=�嘳�d��)
ʶN`<M�N�S .�C�>����	Q��۹Y�<�|^++|�r5��偠�ԗI8�!z'��ֽh�w�م���/����6�ĭ���V#�rٮ��ʘ��lR���2G�q�{D��\������=��T�Փd�u�s��540_Mh��>!��sX�96}�zf��eT[^�1�d\!umiW��i���bݎ|,,?�-u��W��ǻ:��hn'��O4��O��L��G�ʪ�j^���jD�O��vmeH~<�u�0:K��h36j�as���={
_�c�1u���'� �29Iz����<�*�/uQ��]�ʼ��z��zN2IX���n�pu|d5�.4��e
��y;�FTY*S];7'F���d8p��1)9�14��yD{�؛;_��Y�R�]x��	6���yvҸ�mG��)X��A�䉼K��<�@N��}��-�	v�u%�v�=r�r���+~��t�+� ��������b����Z��Q+����5�*��W�1��Vw���?	ƍ��s����� �H����o��Ƴ߸��!�ć�t_u�jտE��8�Z5R]x-���w-�N����d�G��>�	���Z �5�75U�����U
Z����1Pi��;2�z�r@"Ɵ��l��0pK����BS~�J%H����׈�R:b��ߪ�V����h�Ƹ��:YP���q�C��L�0W�}C��dV8����5�+��RFSF�/����bմ�
��}��̨�pֱ���+E�Umn���R�iN6~d%RÌ1�EǆH�-�ָ-a�~��VY�[[�D!jG	��Rr��+!���1?.�=�l�|�	�D҈k�j��6��	��OSc���]�dqq�:���仍��S�h�z��rO�$�(6����;�ĸh�7�@\9_Y�����M���)���'l�	L�Iϝ�s� >*�[z�EP 5����/�nH�%}l��zCvR�����Z�L6&Y�&��	i��Y��``��3�˖Pc&�\���xQ���˴/ƨ| ��l1̔D�%����z�'���`AC����3���#�;�ߧ5`#%��-x��Y	�a�k���ݧԳe.,r�������@q!�KR!ю�Oh���b��̇v�������0k�h�e�n�f���[q�#����)N�Q\}t����M�<?�x�[t�8ҿ�_�}GU���S�Kh�� ��3��x�3��7ŷ��3�R�A2Q�\+�K�l6l�V4�WZM��p�2e��@]f!s�	F�ڜ ��3�ufn��pF�-����z�wz�'D�4>��޸��tAI�V�}��_fX�4	�%�i{]��G��h�WݲV�#��{��D�'�:�0
��+��M�#kz42��6��(�x�Z�j�1�Y�� �C��*a��'Z��2â���PR ���Sx����U�,�ԍ�k�񬧖I�y�q"l��4-rsM��Tp�(,�#�2l,�F'�S�[���ϜێA.��J���/ +_�gp���%Y��[�~zۣy� ����	����%��,�a-�]s�%�}�aSf����M����վFH�2�%��O� _�RT��m�Bvԉ�1�{g��7� /5�s�m�[v�U�������9�ӑ��H�s���F�I��l0(�+4ƙ��m�1�J6�Z͝��b��餑^M��y'�J�2�6�ɳnŐ���w+`�ʷ��)�y�Mr���~�օT�\EߊG���x�'��}�v���&��Sƶ�
�Ƃ�/^�Gb��[�:M�l5σ\ݨ�Eo�O����z��{^*��w+���g�y�ŕ��[�ĭb��4��2�#Q^1�I�5��@���Ri�B�����ũX0�ϊ�W�@��q�a��CWv����wC�YFZa`���A���Vƾ	>z�S��%��X�ҵ��r�&�S�,��2�6�癟0�o���8��V[8��Y���V�]sxS[NYw좟��8�Bz2�Sl�H���h�a����j7�b��WY���k������K��Y.V��ǉԞ!�l��%��X�U$&��t����i���kMj��2�]�`���#��W�5;�Na���^�߾�i���m ɺ��=[�C��#�ǣK)[�H�'i������;�B+ �ϽF��s*o؝�2�B�F��L	ϨR|0����ݯ��q`)���b�F�P��CgR���v�E[䇠��=�迁�p�R|���5;v|����'��̗������
^sS�)PL�����ͣ�^�g~	���c.7�$���򛎐l�������@�C_�������y��h��a>�qU���-j_���Yx�-H�[,I���]O&�m���Sξ���
��y�EP�����c�q�Wm��1�E&��ߩ����I��iK�L9�q�>[�类� w�JUWv�;L�P��j���%�dyp (9�d�V��e:V�VJc��0"�TqK����!ݿ���1 �`c0JX��o�)�y;��Ky�7�e��m�5�xa�KM�0��6��ؚ�{9��mN1�����yD�j�&��@�q�h*4�<��Q9����T����A��!�+r\?�<���`�����9�:���~�W���~������o��}�q�w� �C��5�
����Xf���'Õtk]�A2	�������HkC��H�([��)��j�D�t�s�����Ct��j�Y��o�|�������T������ ��N��S]2�lF~5�=��tv�Zk�ۙ~� �{�X!����U~�6D"Y�.Q�޺�ax�^ŭJ"��s���\kE��ގū=mtw�����l߰%s(�e����;5nճ5_�\l�Hf�)�)ƸQNS��Υ�?�c!���"���ϑ�r��c:5��`�{�L@�>���Z/|�^��QHN��}�������ઉy�^.E���"�{'1ݶ���T�;�Z�9fU�X�*�B���s����N�=ԑV�K��W�3��cs�1��Q���9!i�QoJEb�_"j� �-*O]?>��?��`�!���_�3&���I'~�ƁMa'Q��2�œm�����Og�	��}�����q�d���$��M��>eO��%Q������E���܀B�������K��K<�{�Ls#�4W�Y�"�8�d�7�7:룏�f��qA;X v� {QDtVC*$���
�C���m汣�U��YVT��vq���8��@�nOd�Û*%��h[��O�f����c���h4�����ȼ�r�z�����H�OY�+��Z$�����JӺ�.�>���2X��ϝ��:bw��ƍr 	Ld��-{�(Tb��c����T- �W���}�����|�����H���eg�r۶W�����k�ڡ���8�3���Wl�cc�0��q��W�a
��j�/���7V�@��LsX� �zL$�"�D��.�RC�'���	�c�ن�^Q�=Ck!� �����d�oВg�M�[�>�_7L��j]�������pK��Z�qw������/�Π.R0�d" Ț=wx���/i��y���qf��?��8=��bo�۩F���MId-WJ���{R'n�%�H`X���yRO_�����^�H%�=�+Aj���HUn����+��5eA`'�3D�T�l/����7cԀr�Y�$�$�� ��#j���PY#74��-������u��@�`�^}��߹���dD�^*kbi�B��Y�Ƴ�zWy�Є��|"*��������.�K�:��i��B�l�����.���y�Kx)�Me�$1�ؚM���2�׶k�Ք��ab�U��X�ϥ-�_ϕ��N���@����Bi�Av�4�d��\�/����sJ�6x���C�@�B��E�t��<e��Kʘ�>$�S����I%��.&`�����4�Ց��k���wl��|��yKOxjIqן@m^M#�u�o:gW���#ā���Oԃ-��)D^���鎵K�Zǈ\)����o�:��C"�A1z�j��TkV�W�i��s����.�ca�	��R|���I!�rUǥ����j���v2���4u�Ve^�;�-|�Ie��TC,@g�?�7�����[w��,�]��|��a#��Y��~��� �,�0�l�|1��ro9�7]�cji��d�:7�[gLcQU�C��f���F��(��u�O�/��������9�y<�*�A�S���vS��ě�`Si��n��=^In��ي1p���W�/�����|}��R��r�fc;��ZJ�\E��!�&�a�����g�暕{�[w����_��a��k�X�e�R���p�[n�s5�o�8�W̿���>!��[%�$����.�Cv{/��l�j��n!1DZ���C<"7�����.�P�ai��bG���/��u�+ȕӗ
�!��]H��r4C��B����y���A�j�>?�Ρ1��9W�z7|^����2� �R?�H���j�g�.:�)�#����;s�s?�z����;�|�5�e"���BH��bM���P�+������9bۻ	p�
N�l��!�p+��u
�ܹT.K�]MS}����tT��tc^�%��(v>�P�*��e9�"FͲ{a��@�"���(wڙ��V�FwS7�f�Ĩ�
)�W�!�~�/س� P�@��I�ħ��Whxv��� ^�0.x��J>����l�^��ڮ����o�F.=[���A2��`���O���uu{f��4L��"\��>^ݚ/#��/�٥�?�<�/�Q���|'����;�bUg%��ɬE�r��)��A�k%��_���w�K��GVۮ�����N��_����v]r�w���R��Ȓ�8^A�x��0,F����27����sJ:o�N�e�,����vi�^J��ӷs�4�c�zyk�ٲzm�H������:���L�M��
V q{��#m��m��A��`��A�D���r
$U�A�����ơ&��6 t�b	�襁K�R0��͑c��4�S1�߬"+���;�f�|�l}��,�\����7�"�b��	k�J�<�ƴ�+�i:�	V���j^*�fTnY�0�j��ᝐe2��I��8�*f�o	��E j| �H5�^�´ҫ|�G������^mj�aP)����1��%c�{mv()���r��rWc�^5�\Z�E�#E�E����N���]zg��!1��q���*!6z�A)v��3����D��&�vM�+� �K���l�0j�Y�dG��|��fSֶ���=��D'�� �
g�h0����#w�HREk:]3�i���d9���'h���s9Ѷz4�e��0�j�7Z���8�I_����ۏ2|%�B'�Ok?tR*�ϬWp_um��4��A�w���UUξ~�| '!�_$=,료}��LA��놟z��:��g���8��sbT�Ȉ�C/���x��Ι�k�E�V
S۵.�� ��`�:e�D7c��n�s �t]���M琋�\?��7d:��<���^���(�1�T�1~��O%��'P�WVm����?Y�3yzz�9n�7��`�rʟ9j�%�P�� ɿ�3�������32�E�~ �������rG�M*^���`a@�k̦��W$F�u��4�'nF#�d8K�k4��~��� I8��]ne_����0.��c�-gV��M�c��"�c+z,�l�؝Z@)k�Zm��Sy���U]3��Y�����I��e�����4�}��A����A�)�N��|&����E�d!��х�kc:h�e�<"���Ԑ����2�{��4�W��6p
�+O���0�!3��r��������j1똋*͉����d	�#N���Z���ƶ��'���舾՜e�Z,.��S�,y�D]�0�=�u-=���% �n�P�G�&584Ff��ӕ�K��{�]�l��g�1�E�4j�~��n,Y�N��e ��n���]�Nl�Nm�4�
�	9j��^�]{��^�J]��G����4p�</䏠�y��,QS�r�˟�K�AEZ�7(��G�+��%�L��E�A��yn
��0��e5W�k�"�^?>ŭԈ�ӛK��2�i�Ӏ���������z|k��ҽ�'�ǚU�]��?��P�Y���Ī��e����S}�Z�όS�>��jo������COI�O���	ל������I��hc��]|0* �zn�"�wfx�3�X_�/�:��-?�H�\�D��a���ڰ�tX!L���*�Ӎ
4{��~K����w̱5<'���u?�eBE$<&L(H;8I���R���|2�t.�R���<Sq��˒����H�z�vZ�`3�*Z�H5�H����'�_(g��\n2t�m�`���>������8�s�����ٸ��t�>�7�7�ד��
�N��)����,��wa����9��5��C�d�6 j��J�j�D����J��b���|�Q�F�W��3�~VI|�PEe�x-�]���`K��h�<-��,
-V�SJF�>ٷ�����
ܒ��YQ#�4����?L�}	�C��mw�1�1���8��W�Qw/_&6`�J��X��� Xbyv��j���&2dK�s�SM@�:d[��j7�n#w��z��Q�k�㢖��c^�w&�.����tu���j�B��*��^�?xRҩ48��kI�aDu���BE%#.!�/�����K��m=Ic��mw9�x@�$ୄ�L*�:٦����9]�gE�\Ě��:�;$��qBUn"�d��۪d?��K&��@!��pw<x�������y"K��������
�����νh�/3l�(�ٌ��9U]�wL���<[�1_�t�1"���#ΣC,���ƍ�M��ZXc��]n�b��b���t�x�]A���9޹΄dh��kșyq����E���-���u1����d�g^���?��C�
�cs/a�O��;�6n$�
���'��/\�;��k]1�֥֛p��{$|:���e*�Uh�(�\g�K�����0��0������"IЭ0׺|沊<AHF~��o7i���� �1� �������T���n�IÑ<�3dV���?�7i]MJ�J�"�!��΋�2�� ���>7].V8I[,X�z,�Lz�dY�� |`��`�\����D����Tu�ڞ��e]�¥m��1:���L�Wm�ნ��Μw	b�r��*q:م�h��~3��X�MY�t+k���M�F,���_��6��M��՞<sݔth��b���H��$���n"�)0�yv��V$�$^���Kz�Ǧ�,�+�e�𘀐D�DɌ�i�GĘV��[Y*��Tr�)�~G�ݴM�f@c,�8�i�2��	U��Mu6v����ϐ%ц�8W���ѓ���6���}[J�P'�����:�u��A��r�w2iZB!�i�N�C��]��_�5���-�k�8�$���+v:^�W��J̝����I'}�:�!�Q3�uhf��:��"�v"~W)����b{5�����k[v���9�ˇ���<��eh��$^������*�3���:�(FC���
 ^��yNlB?39�t�G�$-��Ä�� �7��۞�	���|��R��n��Ij)i���ӫE��*�VK����nB�x���3�G�@�|[���������;����:�α��H�~�d��Hm���g�kb"�9��&�Ί������j)���qZ2h�1OwGX�F1�T���M_��,�E�,�$!�1x�#/w��cp�0�2�!���Na�Gq�[��������+�Ɋ���^�T$n )������u�ٙ�1�EFԱ��t�R���?X4Y�_��T��j�"M�MD'�k��٠��#04y�m���h!H��N�+�䥕Q�)���F�T2$�D,�B�%�G�iI��ｍ3sb����<��e�_rَ�K&�J=�gė��H��/k��O4��rx����)^q=h��-pM��A����U�ͩ �	�X������xgW4K��JyYXIR��5ڄ밞����t �0\CB�?9����Ny���TZm���|��]?�
�Ʀ:|��}8e�I�z腳
��	�����/� �O�J�kź�gq���L�=3�+�Ԧ��ϕ�w'4Үji�L�zl)����'a?V��-��-]�H�K��]��G~:/^I����S�Pw�p"�5�<�����}�ɳ��c"�{0}�ۿ�h������h6����<���#� OV�y]y���:�;�H�U2U�2$��:��Ӯi�,X���_F�>�E.�M~���l�f��3�DشY�e�]�ݝu��oR���?7;,�Y��?M$X^��;����X	 ł/�x|7��sH����B����M�އ� /drD4�f���sGA�H�q����|2�����,Gj�(>���댾���`����}s�<�QYR���Ĉ�~�A\:�k������}���D��r�@��;4���w|�+)�XE譆?A��E�h�T���]i?v�p���{��
��T�;F�Ҍ�D&�z�4Dz�m˺���
�������D0B%�e#�Q���O�"#��˞6���!�'�5O��^�<r^_J����`�ƥ�ă����0>�W,�c�� �3�.Y��٘hF����W�9"�ݾ�QVI��E�lbؔ�ēlP"K���$3�\4U]r+:�"���s�d��)Z��Sך�ʸ̖|y�0,��;rl&�'潑L��>��~���{#�DcϽ�P��O5�d���0�Fh�0�~�X��|t=�J��îR
`��L贱L,�Y���r�MĞ��6��(��A[��ߡ���(C���?D����Od�r�*�(5���%	tU�XY9���Q0 �,�f��p+��e0����XξOa@���:��O��:�Iw;��?n�B�������;������A���Mp�gv�d4.܈A���ҭ�u��{~�u���o�,Mw7 ���\/�<ЊpU����(��Y�S$�r��.墒�Ӷ-�׮t������ĘA	��N-^�>�b����O�8$T.ެ��mh�R�a)V��R��&^A�9��t�w�*��Ԭ>�g�Fϴ��@z(�(f
)-ڱU�`;+�^s����wiJ�L��ȑt��$L��B��W��(֛[5w�p��k�{"��V>�}Uo�~5�-�����zư5���d䆊K�_�V��jS�Z��O�xTrU4ħ��3��$�TS2G6��!Е�:;�§�CL~��e���ą���M#��A�q:z�{��H���u���	���3N�
��R�jΥ�;�Î����U�C���N/�`��w����Y�j#c�ڛᙓRc���IH=4�,,���n}��
,N��%L���(Y�vo�㿐���I���ڲ%��q0~���}�D�����]������;���Z<�G�����8�JLo<�ξqF,�,"��:1u��i�;����+q�gY��бa���P��Hh���_�%􈪗szpC�E'=(�C7N�E���v]��ٺ_���?�c�����K$k�7���J��G'V�'~�f������A*+�y���.�8x�}�+��,*�t��A��8�?2�G�?�����e���f1n��*~g�H+�]npd|P����J�#�QU�Ȓz�`
z�
n��[��FPf������i���d��Jg���w�������|qZÿV��nf�0�H��}� Qf�44�}��ف`�Cm@T���+K-<���a��i��)U��Y7RɌת��.DZ\5slɭ���f0�����E�=�lK�AN�/N50|��/,{�wSS�\����v��f�ٓ�,������=���b8���O�f�!'
�b�T,�pj�x�Z�I���w� �E�Ȋ��_Y6(�qD,���d�Ē��6�:��N�� ��<�z�92{�Y��MH!�s���\p�������	����C��׋��b�E|V�0���H�H|<��������{o��G)�#ȟ]}l`%��Q���t2
v��&�IJ�_��s?��ڡ�MR��Qo��w ��H/�B=�&�j/>DNWq������ o���1M��/@�G��w���'��J:��I��рc�[�唔�v�
Y�����V	#(r��RK�[{��E�ђ�V7"�@MBR�lQn����i7�
F�w���(�9W%8�E�b�W	X����9�rø�>ƕ�B6v�[}ꄜ��Gc��k�!�(5�vd.cے�	�g"�Y��@<,-W��X#�I��i���L��D��e%,�>\��~�2�vr8��O����Í���O|��KD��S�7�N�P�N냹jZ8hoEj}q{�	�.6ʭ`�U�B�r���0W�w�%·1����g��d�x��8��z�x�f�ʹe�Ҽ�bp�L��,�n��fyN=�gl_�_��A��x�@�\7�����!忽@ev�ؽL�G��ơ%�C����)�ٹ�{�\�=Դ��gR.Jmf�'�:ş{�e�s3���gLwb�?%�����2�J6l0��1wpq=��2�o7�"�ڤDC0Y��8��Pj���������'�M��'&�����aKo�o�!a�$��U�<���,<s�h����J��M��t�`0�J�Q���*�+#iώ$�_���BE�K�.{����[�&ɘ`(3p�2KMh1��� */��	��}�0\�Ffq~���ǿ6��wmF9�Y��Sb�r�*�K짦�<�yq���W�7	ۅb�g��SM���?�h1�j�/��[��`��,��"b�s���fxv��z9g&%I�ɩ+�_':Q�m�����,��]�^��/�[�`�8C.\n��È �Q���^��E�BC<[n�ɕw�B����H���Ƨ8g��DP��Q9�`ק�!تef�\�0i-Z�#�ZK�'t;G�`t�q3p�����n�ku�:Rr�N�z��)������m��u����/�P%[O����o/��i0�o�ǁ�O`Q~��¬���w�G��=�}`а.���L�m��q���O��s<$y�J�,����~"p��L8��t�UĴ��瑗ǂ"�?n���:~�h;>ڶ�x�*�Lq!deu��^;��|�zN�ۊ�P�$(��J�W��WMC�A��A!���n�fbT�'�5����F�'�aǰ��R+Ӧf���\��J�u��4*�ms_��N^vǔ��Bfg)����X�u ~yH�$���FcE��w�ib̕g�[�R��T[�"bv8��<��R?B�E��
�v:���/=[i��N��U��lN4��V�%ac�j��
��	���-��En9�]z�����LR��0�1�H�%�R�bC7�=��:�(2�q�a�X�&K��1UU�z#�\G9ǸL�Kt?&	�>#{�v���I�c�v�8�Sb��3`�,\È��!l�U����0�UY��T��Ƞ1�*��;k%&�w�A�wz�����k`�h�������O����s�_��1L�y~�Q�	N�E2���<�|3{�
��*k'$W�	IwQR%�E��l)o�C>��i�8���qdƹ-4���kZ�����ʋ$��ڣD�RA��
�ɥ���AV�v��2b���f�5��zQ��l~��5O�2�Y�y�Y�l���ܛ���0Z]�ӵ)Ac��]��C�͞��9��?�p�J~h،ҵ5�6҂a�|QcGB��P1��P��Vw��G��-�7=]P��W��	���� �,!�9�jۨ¢��sve9Oj)K��:�#w�1�Er��ҩF�	�#l�p\����zaUf���_ss����!Z��ܫ��__+"*�@���ub�eMn"��+���@Y�-d@������=>g����Rg.U��̍C�\	_$7�Ro���?��n��M1yp�S�.��bK��`�9����Wv%潾ܐ��)ȅ�G΄�/p#�~�xo'prZ���e/T�L��2��4��p�*|#�%��6������1�q%]��85�K��g���.�%�[n�z4��rL�&@A�h �Ct����L��T�b�c�	S�y�g��ݑ|��}6��pR�Y�@��m������8o�����o�"�W��l���(�.�^��v�������\�ic��1b|��0�?5?��ȯ��x�_H'�b�˚"3��gS_3T�-y��e>B���x+^%���¢&��D����g���1PRq� ���T�h����Q���m�+�dJ���JG��-��]���{��bʸ�����/���.U�_�5;h�D?]�@뜻��좗�O33���ur����Q�o)Zu���2�,� +_� ϥ9o�te�[�o�B؂y�[��UE>��i_�\8��-c%�V�a��_��6�2�Y�a��9�H�PRU4����z܆����x�ʗ��_3!s:m ���}�L�Ƕ������X��"ALV���afG�s.��lu��a"���4W��q��x��R>8�.��'�.d�=���ދ8�x8"GPrl�5������&����b�HXUPfԧ	�
q�GD��j�Ec@�2�X�z��� �(�K�����|�h��1�yX~�<���]�zd׋X�\�ȱ:�?��i,T�{/w��Y��Y�ͣܯY�rG���"�~QZ�Lֹ&J��z����G�������@��L\ɖ*���2ɒ=��u\�7g{���$Fƥ�ҁ���5�%��PY&n�r���� �fn8� ϗ� ��6�H�g�'��Q�;)���s�1T��K�L����ӈ<�R��#Zǿ�|�<uG� +L�^Ԙ��؃�j#��d(��JN�� �ED����Cd8�
���,Q���Hƹ������wpF�=b�����Z�J<��{ghJ����� ��S�8�qe���NT���c�OT��I�>L*�wM��Yz���WgT�?R��Lnf�zjx8ȶ��r$9'+Rا՜�7)��Ny]<!UK��CtE��#���n���8�����ANXk���&��ʵ��n1~�;�#F�w���A�ۂ[�#�Tfm�J�<w�.����q����A�9��y;��]�����L"�X�Khc����,�i�� if�ꚶ<xʂ~oc�6;�ꡰM(�}�N	�k���wg=��pw���w1E\�� ���߻��h��3�X����#F
�O���|�-n����U��/w����K�
MÏ3ȕ�>b����=��i|q��Ӳ;��/�EE���H��nv:��ϱC {�����A��OEE+�шJr����E�����ă�`OL�9Ĳ�RD�A�+��I2�(@�O����؄��a��t@�E�+��J��f���4sΕs�g0h�Ri
P������Q�67���B�K�ݭO�]f���z/�\++���hX������~���G�&�d��d�a9/Dj ��4�h*Q�0����It�K@���39�5ᵉ��ٛa��A�� ��[J������5;Tރ9lʩK����gB��+�(��A�Հ!*��[�-����}E`��O�9�f0�8\)<X����G���pj`�[3�׵u���KǋF���<�aL�7#??�%d�	hM�G��#͠���ǭ�e��T�Sei��4���.�U�v�N�$����?��	(���c~��A�f�<�|X$KhH:�Y�Ꝍ������W�i��.ѡi�s��